778812d46aece3ed3c8e10eebee4bb ����   4 �  org/json/CDL  java/lang/Object <init> ()V Code
  	   LineNumberTable LocalVariableTable this Lorg/json/CDL; getValue *(Lorg/json/JSONTokener;)Ljava/lang/String; 
Exceptions  org/json/JSONException
    org/json/JSONTokener   next ()C  java/lang/StringBuffer
  	  java/lang/StringBuilder  Missing close quote '
  !  " (Ljava/lang/String;)V
  $ % & append (C)Ljava/lang/StringBuilder; ( '.
  * % + -(Ljava/lang/String;)Ljava/lang/StringBuilder;
  - . / toString ()Ljava/lang/String;
  1 2 3 syntaxError ,(Ljava/lang/String;)Lorg/json/JSONException;
  5 % 6 (C)Ljava/lang/StringBuffer;
  -
  9 :  back <  
  > ? @ nextTo (C)Ljava/lang/String; x Lorg/json/JSONTokener; c C q sb Ljava/lang/StringBuffer; StackMapTable MethodParameters rowToJSONArray ,(Lorg/json/JSONTokener;)Lorg/json/JSONArray; M org/json/JSONArray
 L 	
  P  
 L R S T length ()I
 V R W java/lang/String
 L Y Z [ put ((Ljava/lang/Object;)Lorg/json/JSONArray; ] Bad character ' _ ' (
  a % b (I)Ljava/lang/StringBuilder; d ). ja Lorg/json/JSONArray; value Ljava/lang/String; rowToJSONObject A(Lorg/json/JSONArray;Lorg/json/JSONTokener;)Lorg/json/JSONObject;
  l J K
 L n o p toJSONObject +(Lorg/json/JSONArray;)Lorg/json/JSONObject; names s org/json/JSONObject rowToString ((Lorg/json/JSONArray;)Ljava/lang/String;
 L w x y opt (I)Ljava/lang/Object;
  -
 V | } ~ indexOf (I)I
 V � � � charAt (I)C
  � % � ,(Ljava/lang/String;)Ljava/lang/StringBuffer; i I object Ljava/lang/Object; string j toJSONArray ((Ljava/lang/String;)Lorg/json/JSONArray;
  !
  � � K
  � � � @(Lorg/json/JSONArray;Lorg/json/JSONTokener;)Lorg/json/JSONArray; <(Lorg/json/JSONArray;Ljava/lang/String;)Lorg/json/JSONArray;
  � i j jo Lorg/json/JSONObject;
 L � � � optJSONObject (I)Lorg/json/JSONObject;
 r � q � ()Lorg/json/JSONArray;
  � t u
 V � � � valueOf &(Ljava/lang/Object;)Ljava/lang/String;
  � . � <(Lorg/json/JSONArray;Lorg/json/JSONArray;)Ljava/lang/String;
 r � � � *(Lorg/json/JSONArray;)Lorg/json/JSONArray; 
SourceFile CDL.java !               /     *� �    
       .             
            H     �*� < ���	����    �          *   "   ,   '   ,   ,   {�=� Y� N*� <� � 6� 
� 	� *� Y�  � #'� )� ,� 0�-� 4W���-� 7�*� 8;�*� 8*,� =�    
   J    <  =  > < @ > C @ D H F M G R H U J e K  M � E � O � Q � R � T � U    *    � A B    � C D  @ M E D  H E F G  H    
 � ;� 	 �  I    A   	 J K          !     ~� LY� NL*� OM*� >,� +� Q� ,� U� ,� �+,� XW,� ��� � 8
� � � +�*� Y\�  � #^� )� `c� )� ,� 0�*� >���    
   F    `  b  c  d  e * f , h 2 j 8 k ; m A n Q o S q f r r q v t { i    *    ~ A B    v e f   q g h   l C D  H    �  L� ! V" I    A   	 i j           g     +� kM,� ,*� m� �    
   
    �  �          q f      A B    e f  H    �  L@ r I   	 q   A   	 t u    �     ƻ Y� L=� �� 
+,� 4W*� vN-� �-� z:� U� {,� {� +
� {� !� {� � {� � "� I+"� 4W� U66� $� 6 � "� 
+� 4W����+"� 4W� 
+� �W�*� Q��V+
� 4W+� 7�    
   ^    �  �  �  �  �  � " � ( � : � N � b � i � p � v �  � � � � � � � � � � � � � � � � �    R    � e f    � F G  
 � � �   � � �  ( � � h  p 5 S �  s + � �    C D  H   ! 	�  
� I  V� � �  I    e   	 � �           6     � Y*� �� ��    
       �         � h   I    �   	 � K           3     	*� k*� ��    
       �        	 A B   I    A   	 � �           A     *� Y+� �� ��    
       �         q f      � h  I   	 q   �   	 � �           �     6*� 
*� Q� �� LY� NM*+� �N-� � ,-� XW���,� Q� �,�    
   .    �  �  �  �  �  � " � ( � + � 2 � 4 �    *    6 q f     6 A B   ! e f    � �  H    �  L�  r�  I   	 q   A   	 . u           �     /*� �L+� &+� �M,� � Y,� �� ��  ,*� �� )� ,��    
       �  � 
 �  �  � - �         / e f    ) � �    q f  H    � - r I    e   	 . �           �     D*� 
*� Q� �� Y� M>�  +� �:� ,*� �� �� �W�+� Q���,� 7�    
   & 	       ! & 4 ?    4    D q f     D e f   / F G   ( � �  !  � �  H    �   I   	 q   e    �    �